// megafunction wizard: %RAM: 1-PORT%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: altsyncram 

// ============================================================
// File Name: dataMemory.v
// Megafunction Name(s):
// 			altsyncram
//
// Simulation Library Files(s):
// 			altera_mf
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 20.1.0 Build 711 06/05/2020 SJ Lite Edition
// ************************************************************


//Copyright (C) 2020  Intel Corporation. All rights reserved.
//Your use of Intel Corporation's design tools, logic functions 
//and other software and tools, and any partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Intel Program License 
//Subscription Agreement, the Intel Quartus Prime License Agreement,
//the Intel FPGA IP License Agreement, or other applicable license
//agreement, including, without limitation, that your use is for
//the sole purpose of programming logic devices manufactured by
//Intel and sold by Intel or its authorized distributors.  Please
//refer to the applicable agreement for further details, at
//https://fpgasoftware.intel.com/eula.


module dataMemory(address,
	clock,
	data,
	rden,
	wren,
	q);

	input	[31:0]  address;
	input	  clock;
	input	[31:0]  data;
	input	  rden;
	input	  wren;
	output reg	[31:0]  q;

	reg [31:0] DM [255:0]; // 256-word memory

    // Initialize memory with incremental values
    integer i;
    initial begin
        for (i = 0; i < 256; i = i + 1) begin
            DM[i] = i;
        end
    end

    always @(posedge clock) begin
        if (wren)
            DM[address] <= data; // Divide by 4 to get the correct word address
    end

    always @(posedge clock) begin
        if (rden)
            q <= DM[address]; // Divide by 4 to get the correct word address
    end

endmodule